// `include "fulladder.v"
module Adder_64( 
    input [63:0] A,
    input [63:0] B,
    output [63:0] S,
    output cout
);

wire [64:0]Di ;
assign Di[0]=1'b0;

genvar i;
generate
    for(i=0;i<64;i=i+1)
    begin
        fulladder FA(A[i],B[i],Di[i],S[i],Di[i+1]);
    end
endgenerate

assign cout = Di[64]; 

endmodule


// time =0 ,
// a   = 0000000000000000000000000000000000000000000000000000000000010111 ,
// b   = 0000000000000000000000000000000000000000000000000000000000100101 ,
// S   = 0000000000000000000000000000000000000000000000000000000000111100 ,
// Cout = 0 
// time =5 ,
// a   = 1111111111111111111111111111111111111111111111111111111111111101 ,
// b   = 0000000000000000000000000000000000000000000000000000000000001000 ,
// S   = 0000000000000000000000000000000000000000000000000000000000000101 ,
// Cout = 1 
// time =10 ,
// a   = 0000000000000000000000000000000000000000000000000000000111110100 ,
// b   = 1111111111111111111111111111111111111111111111111111111111100111 ,
// S   = 0000000000000000000000000000000000000000000000000000000111011011 ,
// Cout = 1 
// time =15 ,
// a   = 1111111111111111111111111111111111111111111111111111111011010100 ,
// b   = 1111111111111111111111111111111111111111111111111111111110111010 ,
// S   = 1111111111111111111111111111111111111111111111111111111010001110 ,
// Cout = 1 
// time =20 ,
// a   = 1000000000000000000000000000000000000000000000000000000000000000 ,
// b   = 1000000000000000000000000000000000000000000000000000000000000000 ,
// S   = 0000000000000000000000000000000000000000000000000000000000000000 ,
// Cout = 1 
// time =25 ,
// a   = 0010000000000000000000000000000000000000000000000000000000000000 ,
// b   = 0010000000000000000000000000000000000000000000000000000000000000 ,
// S   = 0100000000000000000000000000000000000000000000000000000000000000 ,
// Cout = 0 