`include "fulladder.v"
`include "TwoToFourDecoder.v"
`include "enable.v"
`include "Adder_64.v"
`include "Subtractor_64.v"
`include "And_64.v"
`include "Xor_64.v"

module alu_64(
    input [1:0] alu_fun,
    input [63:0] A,
    input [63:0] B,
    output reg [63:0] valE,
    output reg [2:0] CC // ZF SF OF 
);

wire [63:0] A_add, B_add, A_sub, B_sub, A_and, B_and, A_xor, B_xor;
wire [63:0] AddResult,SubResult, AndResult, XorResult;
wire [3:0] Select;
wire add_cout, sub_cout; 

// 2-to-4 Decoder
TwoToFourDecoder Decoder (
    .A0(alu_fun[0]),
    .A1(alu_fun[1]),
    .D0(Select[0]),
    .D1(Select[1]),
    .D2(Select[2]),
    .D3(Select[3])
);

// Enable Block for Addition
enable EnableAdd (
    .E(Select[0]),
    .A(A),
    .B(B),
    .C(A_add),
    .D(B_add)
);

// Enable Block for Subtraction
enable EnableSub (
    .E(Select[1]),
    .A(A),
    .B(B),
    .C(A_sub),
    .D(B_sub)
);

// Enable Block for AND operation
enable EnableAnd (
    .E(Select[2]),
    .A(A),
    .B(B),
    .C(A_and),
    .D(B_and)
);

// Enable Block for XOR operation
enable EnableXor (
    .E(Select[3]),
    .A(A),
    .B(B),
    .C(A_xor),
    .D(B_xor)
);

// Adder/Subtractor for addition
Adder_64 add (
    .A(A_add),
    .B(B_add),
    .S(AddResult),
    .cout(add_cout) 
);

// Adder/Subtractor for subtraction
Subtractor_64 subtract (
    .A(A_sub),
    .B(B_sub),
    .S(SubResult),
    .cout(sub_cout) 
);

// AND Block
And_64 and1 (
    .A(A_and),
    .B(B_and),
    .AND(AndResult)
);

// XOR Block
Xor_64 xor1 (
    .Out(XorResult),
    .A(A_xor),
    .B(B_xor)
);

//  for selecting the output based on the control signal
always @* begin
    case (alu_fun)
        2'b00: valE = AddResult; 
        2'b01: valE = SubResult;  
        2'b10: valE = AndResult;     
        2'b11: valE = XorResult;     
        default: valE = 64'h0000_0000_0000_0000; 
    endcase
end

always @* begin
    // OF (Over Flow Flag)
   CC[0]=add_cout;
    // SF
    CC[1] = valE[63];
    // ZF (Zero Flag)
    CC[2] = (valE == 64'h0000_0000_0000_0000);
end


endmodule



// time = 0 ,
// alu_fun = 00,
// a   = 0000000000000000000000000000000000000000000000000000000000010111 ,
// b   = 0000000000000000000000000000000000000000000000000000000000100101 ,
// out = 0000000000000000000000000000000000000000000000000000000000111100
// time = 5 ,
// alu_fun = 00,
// a   = 1111111111111111111111111111111111111111111111111111111111111101 ,
// b   = 0000000000000000000000000000000000000000000000000000000000001000 ,
// out = 0000000000000000000000000000000000000000000000000000000000000101
// time = 10 ,
// alu_fun = 00,
// a   = 0000000000000000000000000000000000000000000000000000000111110100 ,
// b   = 1111111111111111111111111111111111111111111111111111111111100111 ,
// out = 0000000000000000000000000000000000000000000000000000000111011011
// time = 15 ,
// alu_fun = 00,
// a   = 1111111111111111111111111111111111111111111111111111111011010100 ,
// b   = 1111111111111111111111111111111111111111111111111111111110111010 ,
// out = 1111111111111111111111111111111111111111111111111111111010001110
// time = 20 ,
// alu_fun = 00,
// a   = 1000000000000000000000000000000000000000000000000000000000000000 ,
// b   = 1000000000000000000000000000000000000000000000000000000000000000 ,
// out = 0000000000000000000000000000000000000000000000000000000000000000
// time = 25 ,
// alu_fun = 00,
// a   = 0010000000000000000000000000000000000000000000000000000000000000 ,
// b   = 0010000000000000000000000000000000000000000000000000000000000000 ,
// out = 0100000000000000000000000000000000000000000000000000000000000000
// time = 30 ,
// alu_fun = 01,
// a   = 0000000000000000000000000000000000000000000000000000000000110110 ,
// b   = 0000000000000000000000000000000000000000000000000000000000101110 ,
// out = 0000000000000000000000000000000000000000000000000000000000001000
// time = 35 ,
// alu_fun = 01,
// a   = 1111111111111111111111111111111111111111111111111111111111111111 ,
// b   = 0000000000000000000000000000000000000000000000000000000000001010 ,
// out = 1111111111111111111111111111111111111111111111111111111111110101
// time = 40 ,
// alu_fun = 01,
// a   = 0000000000000000000000000000000000000000000000000000001111101000 ,
// b   = 1111111111111111111111111111111111111111111111111111111111110001 ,
// out = 0000000000000000000000000000000000000000000000000000001111110111
// time = 45 ,
// alu_fun = 01,
// a   = 1111111111111111111111111111111111111111111111111111111000111001 ,
// b   = 1111111111111111111111111111111111111111111111111111111111010011 ,
// out = 1111111111111111111111111111111111111111111111111111111001100110
// time = 50 ,
// alu_fun = 01,
// a   = 1000000000000000000000000000000000000000000000000000000000000000 ,
// b   = 0100000000000000000000000000000000000000000000000000000000000000 ,
// out = 0100000000000000000000000000000000000000000000000000000000000000
// time = 55 ,
// alu_fun = 01,
// a   = 0100000000000000000000000000000000000000000000000000000000000000 ,
// b   = 1100000000000000000000000000000000000000000000000000000000000000 ,
// out = 1000000000000000000000000000000000000000000000000000000000000000
// time = 60 ,
// alu_fun = 01,
// a   = 0000000000000000000000000000000000000000000000000000000000110110 ,
// b   = 0000000000000000000000000000000000000000000000000000000000110110 ,
// out = 0000000000000000000000000000000000000000000000000000000000000000
// time = 65 ,
// alu_fun = 10,
// a   = 1111111111111111111111111111111111111111111111111111111111111111 ,
// b   = 1111111111111111111111111111111111111111111111111111111111111111 ,
// out = 1111111111111111111111111111111111111111111111111111111111111111
// time = 70 ,
// alu_fun = 10,
// a   = 1111111111111111111111111111111111111111111111111111111111111111 ,
// b   = 0000000000000000000000000000000000000000000000000000000000000000 ,
// out = 0000000000000000000000000000000000000000000000000000000000000000
// time = 75 ,
// alu_fun = 10,
// a   = 1111000011110000111100001111000011110000111100001111000011110000 ,
// b   = 0111100001111000011110000111100001111000011110000111100001111000 ,
// out = 0111000001110000011100000111000001110000011100000111000001110000
// time = 80 ,
// alu_fun = 10,
// a   = 0000000000000000000000000000000000111010110111100110100010110001 ,
// b   = 0000000000000000000000000000000000000111010110111100110100010101 ,
// out = 0000000000000000000000000000000000000010010110100100100000010001
// time = 85 ,
// alu_fun = 10,
// a   = 0000000000000000000000000000000000000111010110111100110100010101 ,
// b   = 1111111111111111111111111111111111000101001000011001011101001111 ,
// out = 0000000000000000000000000000000000000101000000011000010100000101
// time = 90 ,
// alu_fun = 10,
// a   = 1111111111111111111111111111111111111000101001000011001011101011 ,
// b   = 1111111111111111111111111111111111000101001000011001011101001111 ,
// out = 1111111111111111111111111111111111000000001000000001001001001011
// time = 95 ,
// alu_fun = 11,
// a   = 1111111111111111111111111111111111111111111111111111111111111111 ,
// b   = 1111111111111111111111111111111111111111111111111111111111111111 ,
// out = 0000000000000000000000000000000000000000000000000000000000000000
// time = 100 ,
// alu_fun = 11,
// a   = 0000010101010101010101010101010101010101010101010101010101010101 ,
// b   = 0000101010101010101010101010101010101010101010101010101010101010 ,
// out = 0000111111111111111111111111111111111111111111111111111111111111
// time = 105 ,
// alu_fun = 11,
// a   = 0000000000000000000000000000000000000000101111110111011110100000 ,
// b   = 0000000000000000000000000000000000000000000011110111001101000001 ,
// out = 0000000000000000000000000000000000000000101100000000010011100001
// time = 110 ,
// alu_fun = 11,
// a   = 0000000000000000000000000000000000000010101110010010010001010111 ,
// b   = 1111111111111111111111111111111111111111010000001000010101000100 ,
// out = 1111111111111111111111111111111111111101111110011010000100010011
// time = 115 ,
// alu_fun = 11,
// a   = 1111111111111111111111111111111111111111111101110111100011111001 ,
// b   = 1111111111111111111111111111111111111100101010011000111011110000 ,
// out = 0000000000000000000000000000000000000011010111101111011000001001